
module clkdriver (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
