// system_t3.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module system_t3 (
		input  wire        clk_clk,                //             clk.clk
		input  wire [3:0]  parallel_port_0_export, // parallel_port_0.export
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire [11:0] sdram_addr,             //           sdram.addr
		output wire [1:0]  sdram_ba,               //                .ba
		output wire        sdram_cas_n,            //                .cas_n
		output wire        sdram_cke,              //                .cke
		output wire        sdram_cs_n,             //                .cs_n
		inout  wire [15:0] sdram_dq,               //                .dq
		output wire [1:0]  sdram_dqm,              //                .dqm
		output wire        sdram_ras_n,            //                .ras_n
		output wire        sdram_we_n,             //                .we_n
		output wire [7:0]  st2vga_video_data,      //          st2vga.video_data
		output wire        st2vga_video_h_sync,    //                .video_h_sync
		output wire        st2vga_video_v_sync     //                .video_v_sync
	);

	wire         sgdma_0_out_valid;                                                       // sgdma_0:out_valid -> st2vga_0:valid
	wire   [7:0] sgdma_0_out_data;                                                        // sgdma_0:out_data -> st2vga_0:data
	wire         sgdma_0_out_ready;                                                       // st2vga_0:ready -> sgdma_0:out_ready
	wire         sgdma_0_out_startofpacket;                                               // sgdma_0:out_startofpacket -> st2vga_0:startofpacket
	wire         sgdma_0_out_endofpacket;                                                 // sgdma_0:out_endofpacket -> st2vga_0:endofpacket
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                       // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                    // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                    // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [23:0] nios2_gen2_0_data_master_address;                                        // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                     // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                           // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                          // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                      // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [7:0] sgdma_0_m_read_readdata;                                                 // mm_interconnect_0:sgdma_0_m_read_readdata -> sgdma_0:m_read_readdata
	wire         sgdma_0_m_read_waitrequest;                                              // mm_interconnect_0:sgdma_0_m_read_waitrequest -> sgdma_0:m_read_waitrequest
	wire  [31:0] sgdma_0_m_read_address;                                                  // sgdma_0:m_read_address -> mm_interconnect_0:sgdma_0_m_read_address
	wire         sgdma_0_m_read_read;                                                     // sgdma_0:m_read_read -> mm_interconnect_0:sgdma_0_m_read_read
	wire         sgdma_0_m_read_readdatavalid;                                            // mm_interconnect_0:sgdma_0_m_read_readdatavalid -> sgdma_0:m_read_readdatavalid
	wire  [31:0] master_0_master_readdata;                                                // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                             // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                                 // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                                    // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                              // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                                           // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                                   // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                               // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] sgdma_0_descriptor_read_readdata;                                        // mm_interconnect_0:sgdma_0_descriptor_read_readdata -> sgdma_0:descriptor_read_readdata
	wire         sgdma_0_descriptor_read_waitrequest;                                     // mm_interconnect_0:sgdma_0_descriptor_read_waitrequest -> sgdma_0:descriptor_read_waitrequest
	wire  [31:0] sgdma_0_descriptor_read_address;                                         // sgdma_0:descriptor_read_address -> mm_interconnect_0:sgdma_0_descriptor_read_address
	wire         sgdma_0_descriptor_read_read;                                            // sgdma_0:descriptor_read_read -> mm_interconnect_0:sgdma_0_descriptor_read_read
	wire         sgdma_0_descriptor_read_readdatavalid;                                   // mm_interconnect_0:sgdma_0_descriptor_read_readdatavalid -> sgdma_0:descriptor_read_readdatavalid
	wire         sgdma_0_descriptor_write_waitrequest;                                    // mm_interconnect_0:sgdma_0_descriptor_write_waitrequest -> sgdma_0:descriptor_write_waitrequest
	wire  [31:0] sgdma_0_descriptor_write_address;                                        // sgdma_0:descriptor_write_address -> mm_interconnect_0:sgdma_0_descriptor_write_address
	wire         sgdma_0_descriptor_write_write;                                          // sgdma_0:descriptor_write_write -> mm_interconnect_0:sgdma_0_descriptor_write_write
	wire  [31:0] sgdma_0_descriptor_write_writedata;                                      // sgdma_0:descriptor_write_writedata -> mm_interconnect_0:sgdma_0_descriptor_write_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                             // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [23:0] nios2_gen2_0_instruction_master_address;                                 // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                    // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                           // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_chipselect; // mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_chipselect -> parallel_port_0:chipselect
	wire  [31:0] mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_readdata;   // parallel_port_0:readdata -> mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_address;    // mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_address -> parallel_port_0:address
	wire         mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_read;       // mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_read -> parallel_port_0:read
	wire   [3:0] mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_byteenable; // mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_byteenable -> parallel_port_0:byteenable
	wire         mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_write;      // mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_write -> parallel_port_0:write
	wire  [31:0] mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_writedata;  // mm_interconnect_0:parallel_port_0_avalon_parallel_port_slave_writedata -> parallel_port_0:writedata
	wire         mm_interconnect_0_sgdma_0_csr_chipselect;                                // mm_interconnect_0:sgdma_0_csr_chipselect -> sgdma_0:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_0_csr_readdata;                                  // sgdma_0:csr_readdata -> mm_interconnect_0:sgdma_0_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_0_csr_address;                                   // mm_interconnect_0:sgdma_0_csr_address -> sgdma_0:csr_address
	wire         mm_interconnect_0_sgdma_0_csr_read;                                      // mm_interconnect_0:sgdma_0_csr_read -> sgdma_0:csr_read
	wire         mm_interconnect_0_sgdma_0_csr_write;                                     // mm_interconnect_0:sgdma_0_csr_write -> sgdma_0:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_0_csr_writedata;                                 // mm_interconnect_0:sgdma_0_csr_writedata -> sgdma_0:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                 // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;              // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                        // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                          // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                           // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                        // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                             // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                         // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                             // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_controller_0_s1_chipselect;                      // mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_0_s1_readdata;                        // sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_sdram_controller_0_s1_waitrequest;                     // sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_controller_0_s1_address;                         // mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	wire         mm_interconnect_0_sdram_controller_0_s1_read;                            // mm_interconnect_0:sdram_controller_0_s1_read -> sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_0_s1_byteenable;                      // mm_interconnect_0:sdram_controller_0_s1_byteenable -> sdram_controller_0:az_be_n
	wire         mm_interconnect_0_sdram_controller_0_s1_readdatavalid;                   // sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_0_s1_write;                           // mm_interconnect_0:sdram_controller_0_s1_write -> sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_0_s1_writedata;                       // mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	wire         irq_mapper_receiver0_irq;                                                // sgdma_0:csr_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                    // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> master_0:clk_reset_reset
	wire         nios2_gen2_0_debug_reset_request_reset;                                  // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         master_0_master_reset_reset;                                             // master_0:master_reset_reset -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, parallel_port_0:reset, rst_translator:in_reset, sdram_controller_0:reset_n, sgdma_0:system_reset_n, st2vga_0:reset_reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                  // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	system_t3_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                        //          clk.clk
		.clk_reset_reset      (rst_controller_reset_out_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),        //       master.address
		.master_readdata      (master_0_master_readdata),       //             .readdata
		.master_read          (master_0_master_read),           //             .read
		.master_write         (master_0_master_write),          //             .write
		.master_writedata     (master_0_master_writedata),      //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),    //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),  //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),     //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)     // master_reset.reset
	);

	system_t3_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	system_t3_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	system_t3_parallel_port_0 parallel_port_0 (
		.clk        (clk_clk),                                                                 //                        clk.clk
		.reset      (rst_controller_001_reset_out_reset),                                      //                      reset.reset
		.address    (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_readdata),   //                           .readdata
		.in_port    (parallel_port_0_export)                                                   //         external_interface.export
	);

	system_t3_sdram_controller_0 sdram_controller_0 (
		.clk            (clk_clk),                                               //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                            //  wire.export
		.zs_ba          (sdram_ba),                                              //      .export
		.zs_cas_n       (sdram_cas_n),                                           //      .export
		.zs_cke         (sdram_cke),                                             //      .export
		.zs_cs_n        (sdram_cs_n),                                            //      .export
		.zs_dq          (sdram_dq),                                              //      .export
		.zs_dqm         (sdram_dqm),                                             //      .export
		.zs_ras_n       (sdram_ras_n),                                           //      .export
		.zs_we_n        (sdram_we_n)                                             //      .export
	);

	system_t3_sgdma_0 sgdma_0 (
		.clk                           (clk_clk),                                  //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),      //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_0_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_0_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_0_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_0_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_0_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_0_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_0_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_0_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_0_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_0_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_0_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_0_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_0_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_0_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_0_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                 //          csr_irq.irq
		.m_read_readdata               (sgdma_0_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_0_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_0_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_0_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_0_m_read_read),                      //                 .read
		.out_data                      (sgdma_0_out_data),                         //              out.data
		.out_valid                     (sgdma_0_out_valid),                        //                 .valid
		.out_ready                     (sgdma_0_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_0_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_0_out_startofpacket)                 //                 .startofpacket
	);

	st2vga #(
		.WIDTH (8),
		.DIV   (4)
	) st2vga_0 (
		.ready         (sgdma_0_out_ready),                   // avalon_streaming_sink.ready
		.valid         (sgdma_0_out_valid),                   //                      .valid
		.data          (sgdma_0_out_data),                    //                      .data
		.startofpacket (sgdma_0_out_startofpacket),           //                      .startofpacket
		.endofpacket   (sgdma_0_out_endofpacket),             //                      .endofpacket
		.reset_reset_n (~rst_controller_001_reset_out_reset), //            reset_sink.reset_n
		.clk_clk       (clk_clk),                             //            clock_sink.clk
		.video_data    (st2vga_video_data),                   //                   vga.video_data
		.video_h_sync  (st2vga_video_h_sync),                 //                      .video_h_sync
		.video_v_sync  (st2vga_video_v_sync)                  //                      .video_v_sync
	);

	system_t3_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                                 //                                  clk_0_clk.clk
		.master_0_clk_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                                      //   master_0_clk_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                                      //   nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.master_0_master_address                               (master_0_master_address),                                                 //                            master_0_master.address
		.master_0_master_waitrequest                           (master_0_master_waitrequest),                                             //                                           .waitrequest
		.master_0_master_byteenable                            (master_0_master_byteenable),                                              //                                           .byteenable
		.master_0_master_read                                  (master_0_master_read),                                                    //                                           .read
		.master_0_master_readdata                              (master_0_master_readdata),                                                //                                           .readdata
		.master_0_master_readdatavalid                         (master_0_master_readdatavalid),                                           //                                           .readdatavalid
		.master_0_master_write                                 (master_0_master_write),                                                   //                                           .write
		.master_0_master_writedata                             (master_0_master_writedata),                                               //                                           .writedata
		.nios2_gen2_0_data_master_address                      (nios2_gen2_0_data_master_address),                                        //                   nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                  (nios2_gen2_0_data_master_waitrequest),                                    //                                           .waitrequest
		.nios2_gen2_0_data_master_byteenable                   (nios2_gen2_0_data_master_byteenable),                                     //                                           .byteenable
		.nios2_gen2_0_data_master_read                         (nios2_gen2_0_data_master_read),                                           //                                           .read
		.nios2_gen2_0_data_master_readdata                     (nios2_gen2_0_data_master_readdata),                                       //                                           .readdata
		.nios2_gen2_0_data_master_write                        (nios2_gen2_0_data_master_write),                                          //                                           .write
		.nios2_gen2_0_data_master_writedata                    (nios2_gen2_0_data_master_writedata),                                      //                                           .writedata
		.nios2_gen2_0_data_master_debugaccess                  (nios2_gen2_0_data_master_debugaccess),                                    //                                           .debugaccess
		.nios2_gen2_0_instruction_master_address               (nios2_gen2_0_instruction_master_address),                                 //            nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest           (nios2_gen2_0_instruction_master_waitrequest),                             //                                           .waitrequest
		.nios2_gen2_0_instruction_master_read                  (nios2_gen2_0_instruction_master_read),                                    //                                           .read
		.nios2_gen2_0_instruction_master_readdata              (nios2_gen2_0_instruction_master_readdata),                                //                                           .readdata
		.nios2_gen2_0_instruction_master_readdatavalid         (nios2_gen2_0_instruction_master_readdatavalid),                           //                                           .readdatavalid
		.sgdma_0_descriptor_read_address                       (sgdma_0_descriptor_read_address),                                         //                    sgdma_0_descriptor_read.address
		.sgdma_0_descriptor_read_waitrequest                   (sgdma_0_descriptor_read_waitrequest),                                     //                                           .waitrequest
		.sgdma_0_descriptor_read_read                          (sgdma_0_descriptor_read_read),                                            //                                           .read
		.sgdma_0_descriptor_read_readdata                      (sgdma_0_descriptor_read_readdata),                                        //                                           .readdata
		.sgdma_0_descriptor_read_readdatavalid                 (sgdma_0_descriptor_read_readdatavalid),                                   //                                           .readdatavalid
		.sgdma_0_descriptor_write_address                      (sgdma_0_descriptor_write_address),                                        //                   sgdma_0_descriptor_write.address
		.sgdma_0_descriptor_write_waitrequest                  (sgdma_0_descriptor_write_waitrequest),                                    //                                           .waitrequest
		.sgdma_0_descriptor_write_write                        (sgdma_0_descriptor_write_write),                                          //                                           .write
		.sgdma_0_descriptor_write_writedata                    (sgdma_0_descriptor_write_writedata),                                      //                                           .writedata
		.sgdma_0_m_read_address                                (sgdma_0_m_read_address),                                                  //                             sgdma_0_m_read.address
		.sgdma_0_m_read_waitrequest                            (sgdma_0_m_read_waitrequest),                                              //                                           .waitrequest
		.sgdma_0_m_read_read                                   (sgdma_0_m_read_read),                                                     //                                           .read
		.sgdma_0_m_read_readdata                               (sgdma_0_m_read_readdata),                                                 //                                           .readdata
		.sgdma_0_m_read_readdatavalid                          (sgdma_0_m_read_readdatavalid),                                            //                                           .readdatavalid
		.nios2_gen2_0_debug_mem_slave_address                  (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                  //               nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                    //                                           .write
		.nios2_gen2_0_debug_mem_slave_read                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                     //                                           .read
		.nios2_gen2_0_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                 //                                           .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                //                                           .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),               //                                           .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),              //                                           .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),              //                                           .debugaccess
		.onchip_memory2_0_s1_address                           (mm_interconnect_0_onchip_memory2_0_s1_address),                           //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                             (mm_interconnect_0_onchip_memory2_0_s1_write),                             //                                           .write
		.onchip_memory2_0_s1_readdata                          (mm_interconnect_0_onchip_memory2_0_s1_readdata),                          //                                           .readdata
		.onchip_memory2_0_s1_writedata                         (mm_interconnect_0_onchip_memory2_0_s1_writedata),                         //                                           .writedata
		.onchip_memory2_0_s1_byteenable                        (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                        //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                        (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                        //                                           .chipselect
		.onchip_memory2_0_s1_clken                             (mm_interconnect_0_onchip_memory2_0_s1_clken),                             //                                           .clken
		.parallel_port_0_avalon_parallel_port_slave_address    (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_address),    // parallel_port_0_avalon_parallel_port_slave.address
		.parallel_port_0_avalon_parallel_port_slave_write      (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_write),      //                                           .write
		.parallel_port_0_avalon_parallel_port_slave_read       (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_read),       //                                           .read
		.parallel_port_0_avalon_parallel_port_slave_readdata   (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_readdata),   //                                           .readdata
		.parallel_port_0_avalon_parallel_port_slave_writedata  (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_writedata),  //                                           .writedata
		.parallel_port_0_avalon_parallel_port_slave_byteenable (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_byteenable), //                                           .byteenable
		.parallel_port_0_avalon_parallel_port_slave_chipselect (mm_interconnect_0_parallel_port_0_avalon_parallel_port_slave_chipselect), //                                           .chipselect
		.sdram_controller_0_s1_address                         (mm_interconnect_0_sdram_controller_0_s1_address),                         //                      sdram_controller_0_s1.address
		.sdram_controller_0_s1_write                           (mm_interconnect_0_sdram_controller_0_s1_write),                           //                                           .write
		.sdram_controller_0_s1_read                            (mm_interconnect_0_sdram_controller_0_s1_read),                            //                                           .read
		.sdram_controller_0_s1_readdata                        (mm_interconnect_0_sdram_controller_0_s1_readdata),                        //                                           .readdata
		.sdram_controller_0_s1_writedata                       (mm_interconnect_0_sdram_controller_0_s1_writedata),                       //                                           .writedata
		.sdram_controller_0_s1_byteenable                      (mm_interconnect_0_sdram_controller_0_s1_byteenable),                      //                                           .byteenable
		.sdram_controller_0_s1_readdatavalid                   (mm_interconnect_0_sdram_controller_0_s1_readdatavalid),                   //                                           .readdatavalid
		.sdram_controller_0_s1_waitrequest                     (mm_interconnect_0_sdram_controller_0_s1_waitrequest),                     //                                           .waitrequest
		.sdram_controller_0_s1_chipselect                      (mm_interconnect_0_sdram_controller_0_s1_chipselect),                      //                                           .chipselect
		.sgdma_0_csr_address                                   (mm_interconnect_0_sgdma_0_csr_address),                                   //                                sgdma_0_csr.address
		.sgdma_0_csr_write                                     (mm_interconnect_0_sgdma_0_csr_write),                                     //                                           .write
		.sgdma_0_csr_read                                      (mm_interconnect_0_sgdma_0_csr_read),                                      //                                           .read
		.sgdma_0_csr_readdata                                  (mm_interconnect_0_sgdma_0_csr_readdata),                                  //                                           .readdata
		.sgdma_0_csr_writedata                                 (mm_interconnect_0_sgdma_0_csr_writedata),                                 //                                           .writedata
		.sgdma_0_csr_chipselect                                (mm_interconnect_0_sgdma_0_csr_chipselect)                                 //                                           .chipselect
	);

	system_t3_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (master_0_master_reset_reset),            // reset_in2.reset
		.clk            (),                                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.reset_in2      (master_0_master_reset_reset),            // reset_in2.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
