
module clkinter (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
